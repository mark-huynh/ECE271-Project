//Test verilog file

//Try editing this and commiting your changes and I can check if your changes came through.
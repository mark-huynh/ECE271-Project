//Test verilog file

//Try editing this and commiting your changes and I can check if your changes came through.

//Hey I added this can you see it?
module decoder (input s,
					output q);
	
	if(s == 1) q = 1;
	
endmodule
module decoder (input logic s, en
					output logic q);
	
//	always@(posedge en)
//	if(s == 1) 
//	q = 1;
//	
endmodule 